`include "my_intf.sv"
`include "my_trans.sv"
`include "my_sequencer.sv"
`include "my_sequence.sv"
`include "my_isr_seq.sv"
`include "my_driver.sv"
`include "my_monitor.sv"
`include "my_agent.sv"
`include "my_scb.sv"
`include "my_env.sv"
`include "my_driver_callback.sv"
`include "drv_print_cb.sv"
`include "my_test.sv"
`include "test_wr_only.sv"
`include "test_rd_only.sv"
`include "test_rd_wr.sv"
`include "test_rd_wr_con.sv"
`include "test_rd_wr_mix.sv"
`include "test_rd_wr_with_cb.sv"
`include "test_rd_wr_with_DPI.sv"
`include "test_full_interrupt.sv"
`include "test_empty_interrupt.sv"
